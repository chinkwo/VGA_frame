module	vga_module(
		input		wire			sclk			,
		input		wire			rst_n			,
		input		wire			vga_clk		,
		input		wire[7:0]	dout			,
		output	reg				h_sync		,
		output	reg				v_sync		,
		output	wire		area		,
		output	reg[2:0]	r					,
		output	reg[2:0]	g					,
		output	reg[1:0]	b
);
//-----------------------------------------------------------//
// ˮƽɨ��������趨1024*768 60Hz VGA
//-----------------------------------------------------------//
//parameter LinePeriod =1344;            //��������
//parameter H_SyncPulse=136;             //��ͬ�����壨Sync a��
//parameter H_BackPorch=160;             //��ʾ���أ�Back porch b��
//parameter H_ActivePix=1024;            //��ʾʱ��Σ�Display interval c��
//parameter H_FrontPorch=24;             //��ʾǰ�أ�Front porch d��
//parameter Hde_start=296;
//parameter Hde_end=1320;

//-----------------------------------------------------------//
// ��ֱɨ��������趨1024*768 60Hz VGA
//-----------------------------------------------------------//
//parameter FramePeriod =806;           //��������
//parameter V_SyncPulse=6;              //��ͬ�����壨Sync o��
//parameter V_BackPorch=29;             //��ʾ���أ�Back porch p��
//parameter V_ActivePix=768;            //��ʾʱ��Σ�Display interval q��
//parameter V_FrontPorch=3;             //��ʾǰ�أ�Front porch r��
//parameter Vde_start=35;
//parameter Vde_end=803;

//-----------------------------------------------------------//
// ˮƽɨ��������趨800*600 VGA
//-----------------------------------------------------------//
//parameter LinePeriod =1056;           //��������
//parameter H_SyncPulse=128;            //��ͬ�����壨Sync a��
//parameter H_BackPorch=88;             //��ʾ���أ�Back porch b��
//parameter H_ActivePix=800;            //��ʾʱ��Σ�Display interval c��
//parameter H_FrontPorch=40;            //��ʾǰ�أ�Front porch d��

//-----------------------------------------------------------//
// ��ֱɨ��������趨800*600 VGA
//-----------------------------------------------------------//
//parameter FramePeriod =628;           //��������
//parameter V_SyncPulse=4;              //��ͬ�����壨Sync o��
//parameter V_BackPorch=23;             //��ʾ���أ�Back porch p��
//parameter V_ActivePix=600;            //��ʾʱ��Σ�Display interval q��
//parameter V_FrontPorch=1;             //��ʾǰ�أ�Front porch r��

//-----------------------------------------------------------//
// ˮƽɨ��������趨640*480 60Hz VGA
//-----------------------------------------------------------//
parameter LinePeriod =800;            //��������
parameter H_SyncPulse=96;             //��ͬ�����壨Sync a��
parameter H_BackPorch=40;             //��ʾ���أ�Back porch b��
parameter H_ActivePix=640;            //��ʾʱ��Σ�Display interval c��
parameter H_FrontPorch=8;             //��ʾǰ�أ�Front porch d��
parameter Hde_start=144;
parameter Hde_end=784;

//-----------------------------------------------------------//
// ��ֱɨ��������趨640*480 60Hz VGA
//-----------------------------------------------------------//
parameter FramePeriod =525;           //��������
parameter V_SyncPulse=2;              //��ͬ�����壨Sync o��
parameter V_BackPorch=25;             //��ʾ���أ�Back porch p��
parameter V_ActivePix=480;            //��ʾʱ��Σ�Display interval q��
parameter V_FrontPorch=2;             //��ʾǰ�أ�Front porch r��
parameter Vde_start=35;
parameter Vde_end=515;
parameter MOVE_SPEED=(FramePeriod*LinePeriod)-1;

	reg[9:0]			h_cnt		;	//h_cnt==LinePeriod
	reg[9:0]			v_cnt		;	//v_cnt==FramePeriod
	wire					area1		;
	wire					area2		;
	wire					area3		;
//H_cnt�м�����	
always@(posedge	vga_clk	or	negedge	rst_n)
		if(rst_n==0)
			h_cnt	<=	1;
		else	if(h_cnt==LinePeriod)
			h_cnt	<=	1;
		else	if(vga_clk==1)
			h_cnt	<=	h_cnt	+	1;
			
			
//V_cnt�м�����				
always@(posedge	vga_clk	or	negedge	rst_n)
		if(rst_n==0)
			v_cnt	<=	1;
		else	if(v_cnt==FramePeriod&&h_cnt==LinePeriod)
			v_cnt	<=	1;
		else	if(h_cnt==LinePeriod)
			v_cnt	<=	v_cnt	+	1;
			
//h_sync��ͬ���ź�
always@(posedge	vga_clk	or	negedge	rst_n)
		if(rst_n==0)
			h_sync	<=	0;
		else	if(h_cnt==1)
			h_sync	<=	1;
		else	if(h_cnt>=H_SyncPulse)
			h_sync	<=	0;
			
//v_sync��ͬ���ź�
always@(posedge	vga_clk	or	negedge	rst_n)
		if(rst_n==0)
			v_sync	<=	0;
		else	if(v_cnt==1)
			v_sync	<=	1;
		else	if(v_cnt==V_SyncPulse)
			v_sync	<=	0;
/********************************************************************/			
/***************************��̬��������*************************/
	reg					flag_x	;
	reg					flag_y	;
	reg[9:0]		X0			;
	reg[9:0]		Y0			;
	reg[30:0]		cnt_move;
	parameter			X=144	;//������ԭ�㶨��
	parameter			Y=35	;//������ԭ�㶨��
	
//flag_x����	
always@(posedge	vga_clk	or	negedge	rst_n)
	if(rst_n==0)
		flag_x	<=	0;
	else	if((X0)==Hde_start)
		flag_x	<=	1;
	else	if((X0+200)==Hde_end)
		flag_x	<=	0;
			
//flag_x����
always@(posedge	vga_clk	or	negedge	rst_n)
	if(rst_n==0)
		flag_y	<=	0;
	else	if((Y0)==Vde_start)
		flag_y	<=	1;
	else	if((Y0+200)==Vde_end)
		flag_y	<=	0;

//X0����
always@(posedge	vga_clk	or	negedge	rst_n)
	if(rst_n==0)
		X0	<=	X;
	else	if(cnt_move==MOVE_SPEED)
		begin	
			if(flag_x==1)
				X0	<=	X0	+	1;
			else	if(flag_x==0)
				X0	<=	X0-1;
		end

//Y0����
always@(posedge	vga_clk	or	negedge	rst_n)
	if(rst_n==0)
		Y0	<=	Y;
	else	if(cnt_move==MOVE_SPEED)
		begin	
			if(flag_y==1) 
				Y0	<=	Y0	+	1;
			else	if(flag_y==0)
				Y0	<=	Y0-1;
		end				

//cnt_move
always@(posedge	vga_clk	or	negedge	rst_n)
if(rst_n==0)
	cnt_move	<=	0;
else	if(cnt_move<MOVE_SPEED)
	cnt_move	<=	cnt_move+1;
else
	cnt_move	<=	0;

      	
		
/********************************************************************/	

//area������
parameter		R1	=	100	;
parameter		R2	=	50	;
assign	area1	=	(((h_cnt-X0)*(h_cnt-X0)+(v_cnt-Y0)*(v_cnt-Y0))<=(R1*R1));
assign	area2	=	((R2*R2)<=((h_cnt-X0)*(h_cnt-X0)+(v_cnt-Y0)*(v_cnt-Y0)));
assign	area	=	((h_cnt-X0<200)&&(v_cnt-Y0<200));
assign	area4	=	((h_cnt-X<200)&&(v_cnt-Y<200));

//rgb��ֵ
always@(posedge	vga_clk	or	negedge	rst_n)
if(rst_n==0)
		{r,g,b}	<=	8'b000_000_00;
//else	if(area1&&area2)
//		{r,g,b}	<=	8'b011_011_01;
else	if(area)
		{r,g,b}	<=	dout; 
else	if(h_cnt>=Hde_start&&h_cnt<=Hde_end&&v_cnt>=Vde_start&&v_cnt<=Vde_start+160)
		{r,g,b}	<=	8'b111_000_00;
else	if(h_cnt>=Hde_start&&h_cnt<=Hde_end&&v_cnt>=Vde_start&&v_cnt<=Vde_start+320)
		{r,g,b}	<=	8'b000_111_000; 
else	if(h_cnt>=Hde_start&&h_cnt<=Hde_end&&v_cnt>=Vde_start&&v_cnt<=Vde_start+480)
		{r,g,b}	<=	8'b000_000_11;
else	
		{r,g,b}	<=	8'b000_000_00;	
	
		
endmodule